module core_top();




endmodule 