module top();

endmodule 