module stage_decode(
    input [31:0] if_pc, // a la memoria rom y a reg de decode
    input [31:0] de_pc, de_pc_plus4
    
);



endmodule